//`define RISCV
`define ZEPHYR
//`define ZEPHYR_SYNC
//`define ZEPHYR_PHIL
//`define TESTN
//`define DHRYSTONE
//`define INT_TEST
//`define PG_TEST

