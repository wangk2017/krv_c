//`define RISCV
`define BREAKPOINT
//`define SINGLE_STEP
//`define EBREAK
//`define DBG_REF
//`define ZEPHYR
//`define ZEPHYR_SYNC
//`define ZEPHYR_PHIL
//`define TESTN
//`define DHRYSTONE
//`define INT_TEST
//`define PG_TEST

